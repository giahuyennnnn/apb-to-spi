package spi_regmodel_pkg;

	import uvm_pkg::*;
	import apb_pkg::*;
	import spi_register_pkg::*;

	`include "spi_reg2apb_adapter.sv"
	`include "spi_reg_block.sv"
endpackage
