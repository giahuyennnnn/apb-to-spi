package spi_register_pkg;

	import uvm_pkg::*;

	`include "spi_LCR_reg.sv"
	`include "spi_DLR_reg.sv"
	`include "spi_IER_reg.sv"
	`include "spi_FSR_reg.sv"
	`include "spi_TBR_reg.sv"
	`include "spi_RBR_reg.sv"
endpackage
