interface spi_if();
   logic       SCLK;
   logic       MOSI;
   logic       MISO;
   logic [3:0] SS;
endinterface
