`ifndef GUARD_SPI_TEST_PKG__SV
`define GUARD_SPI_TEST_PKG__SV

package test_pkg;
	import uvm_pkg::*;
	import apb_pkg::*;
	import env_pkg::*;
	import seq_pkg::*;
	import spi_regmodel_pkg::*;
	import spi_pkg::*;

	`include "spi_base_test.sv"

   `include "reg_default_test.sv"
   `include "reg_rw_test.sv"
   `include "reg_rsvd_test.sv"

	`include "spi_non_8bit_cpol0_cpha0_slave0_test.sv"
	`include "spi_non_8bit_cpol0_cpha0_slave1_test.sv"
	`include "spi_non_8bit_cpol0_cpha0_slave2_test.sv"
	`include "spi_non_8bit_cpol0_cpha0_slave3_test.sv"
	`include "spi_non_8bit_cpol0_cpha1_slave0_test.sv"
	`include "spi_non_8bit_cpol0_cpha1_slave1_test.sv"
	`include "spi_non_8bit_cpol0_cpha1_slave2_test.sv"
	`include "spi_non_8bit_cpol0_cpha1_slave3_test.sv"
	`include "spi_non_8bit_cpol1_cpha0_slave0_test.sv"
	`include "spi_non_8bit_cpol1_cpha0_slave1_test.sv"
	`include "spi_non_8bit_cpol1_cpha0_slave2_test.sv"
	`include "spi_non_8bit_cpol1_cpha0_slave3_test.sv"
	`include "spi_non_8bit_cpol1_cpha1_slave0_test.sv"
	`include "spi_non_8bit_cpol1_cpha1_slave1_test.sv"
	`include "spi_non_8bit_cpol1_cpha1_slave2_test.sv"
	`include "spi_non_8bit_cpol1_cpha1_slave3_test.sv"
	`include "spi_non_16bit_cpol0_cpha0_slave0_test.sv"
	`include "spi_non_16bit_cpol0_cpha0_slave1_test.sv"
	`include "spi_non_16bit_cpol0_cpha0_slave2_test.sv"
	`include "spi_non_16bit_cpol0_cpha0_slave3_test.sv"
	`include "spi_non_16bit_cpol0_cpha1_slave0_test.sv"
	`include "spi_non_16bit_cpol0_cpha1_slave1_test.sv"
	`include "spi_non_16bit_cpol0_cpha1_slave2_test.sv"
	`include "spi_non_16bit_cpol0_cpha1_slave3_test.sv"
	`include "spi_non_16bit_cpol1_cpha0_slave0_test.sv"
	`include "spi_non_16bit_cpol1_cpha0_slave1_test.sv"
	`include "spi_non_16bit_cpol1_cpha0_slave2_test.sv"
	`include "spi_non_16bit_cpol1_cpha0_slave3_test.sv"
	`include "spi_non_16bit_cpol1_cpha1_slave0_test.sv"
	`include "spi_non_16bit_cpol1_cpha1_slave1_test.sv"
	`include "spi_non_16bit_cpol1_cpha1_slave2_test.sv"
	`include "spi_non_16bit_cpol1_cpha1_slave3_test.sv"
	`include "spi_en_8bit_cpol0_cpha0_slave0_test.sv"
	`include "spi_en_8bit_cpol0_cpha0_slave1_test.sv"
	`include "spi_en_8bit_cpol0_cpha0_slave2_test.sv"
	`include "spi_en_8bit_cpol0_cpha0_slave3_test.sv"
	`include "spi_en_8bit_cpol0_cpha1_slave0_test.sv"
	`include "spi_en_8bit_cpol0_cpha1_slave1_test.sv"
	`include "spi_en_8bit_cpol0_cpha1_slave2_test.sv"
	`include "spi_en_8bit_cpol0_cpha1_slave3_test.sv"
	`include "spi_en_8bit_cpol1_cpha0_slave0_test.sv"
	`include "spi_en_8bit_cpol1_cpha0_slave1_test.sv"
	`include "spi_en_8bit_cpol1_cpha0_slave2_test.sv"
	`include "spi_en_8bit_cpol1_cpha0_slave3_test.sv"
	`include "spi_en_8bit_cpol1_cpha1_slave0_test.sv"
	`include "spi_en_8bit_cpol1_cpha1_slave1_test.sv"
	`include "spi_en_8bit_cpol1_cpha1_slave2_test.sv"
	`include "spi_en_8bit_cpol1_cpha1_slave3_test.sv"
	`include "spi_en_16bit_cpol0_cpha0_slave0_test.sv"
	`include "spi_en_16bit_cpol0_cpha0_slave1_test.sv"
	`include "spi_en_16bit_cpol0_cpha0_slave2_test.sv"
	`include "spi_en_16bit_cpol0_cpha0_slave3_test.sv"
	`include "spi_en_16bit_cpol0_cpha1_slave0_test.sv"
	`include "spi_en_16bit_cpol0_cpha1_slave1_test.sv"
	`include "spi_en_16bit_cpol0_cpha1_slave2_test.sv"
	`include "spi_en_16bit_cpol0_cpha1_slave3_test.sv"
	`include "spi_en_16bit_cpol1_cpha0_slave0_test.sv"
	`include "spi_en_16bit_cpol1_cpha0_slave1_test.sv"
	`include "spi_en_16bit_cpol1_cpha0_slave2_test.sv"
	`include "spi_en_16bit_cpol1_cpha0_slave3_test.sv"
	`include "spi_en_16bit_cpol1_cpha1_slave0_test.sv"
	`include "spi_en_16bit_cpol1_cpha1_slave1_test.sv"
	`include "spi_en_16bit_cpol1_cpha1_slave2_test.sv"
	`include "spi_en_16bit_cpol1_cpha1_slave3_test.sv"
	
	`include "interrupt_rx_full_en_test.sv"
	`include "interrupt_rx_full_dis_test.sv"
	`include "interrupt_rx_empty_en_test.sv"
	`include "interrupt_rx_empty_dis_test.sv"
	`include "interrupt_tx_full_en_test.sv"
	`include "interrupt_tx_full_dis_test.sv"
	`include "interrupt_tx_empty_en_test.sv"
	`include "interrupt_tx_empty_dis_test.sv"
	
	`include "APB_20MHz_test.sv"
	`include "APB_50MHz_test.sv"
	`include "APB_100MHz_test.sv"
	`include "APB_random_test.sv"
	
	`include "dynamic_config_test.sv"
	`include "mismatch_word_test.sv"
	`include "mismatch_cpol_test.sv"
	`include "mismatch_cpha_test.sv"
	`include "mismatch_slave_test.sv"
	
	`include "spi_busy_cfg_LCR_test.sv"
	`include "spi_busy_cfg_DLR_test.sv"
endpackage
`endif
